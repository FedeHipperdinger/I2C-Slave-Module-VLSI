*** SPICE deck for cell XOR{sch} from library ADCD_Hipperdinger
*** Created on mié may. 22, 2024 16:19:23
*** Last revised on mié may. 22, 2024 20:35:43
*** Written on mié may. 22, 2024 20:35:46 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include C:\Users\feder\Desktop\UNS\5to_anio\2do_cuatrimestre\ADCD\Electric\Electric_libs\Modelos_Transistores.txt

*** SUBCIRCUIT ADCD_Hipperdinger__NAND FROM CELL NAND{sch}
.SUBCKT ADCD_Hipperdinger__NAND gnd Va Vb vdd Vout
** GLOBAL gnd
** GLOBAL vdd
Mnmos-4@0 Vout Vb net@3 net@3 NMOS L=0.6U W=1.8U
Mnmos-4@1 net@3 Va gnd gnd NMOS L=0.6U W=1.8U
Mpmos-4@0 vdd Vb Vout vdd PMOS L=0.6U W=3U
Mpmos-4@1 vdd Va Vout pmos-4@1_b PMOS L=0.6U W=3U

* Spice Code nodes in cell cell 'NAND{sch}'
#.INCLUDE Modelos_Transistores.txt
#.PARAM SUPPLY=5v
#VDD VDD 0 DC 'SUPPLY'
#Va Va 0 PULSE 0 'SUPPLY' 100MS 10MS 10MS 200MS 500MS
#Vb Vb 0 PULSE 0 'SUPPLY' 150MS 10MS 10MS 200MS 500MS
#.TRAN 1MS 600MS
.ENDS ADCD_Hipperdinger__NAND

.global gnd vdd

*** TOP LEVEL CELL: XOR{sch}
XNAND@0 gnd net@8 net@5 vdd Vout ADCD_Hipperdinger__NAND
XNAND@1 gnd Va net@0 vdd net@8 ADCD_Hipperdinger__NAND
XNAND@2 gnd net@0 Vb vdd net@5 ADCD_Hipperdinger__NAND
XNAND@3 gnd Va Vb vdd net@0 ADCD_Hipperdinger__NAND
.END
