*** SPICE deck for cell 3b_counter{sch} from library ADCD_Hipperdinger
*** Created on mar jun. 25, 2024 20:47:21
*** Last revised on mar jun. 25, 2024 23:20:23
*** Written on mar jun. 25, 2024 23:20:30 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include C:\Users\feder\Desktop\UNS\5to_anio\2do_cuatrimestre\ADCD\Electric\Electric_libs\Modelos_Transistores.txt

*** SUBCIRCUIT ADCD_Hipperdinger__inv FROM CELL inv{sch}
.SUBCKT ADCD_Hipperdinger__inv gnd vdd Vin Vout
** GLOBAL gnd
** GLOBAL vdd
Mnmos-4@0 Vout Vin gnd gnd NMOS L=0.6U W=1.8U
Mpmos-4@0 vdd Vin Vout vdd PMOS L=0.6U W=3U

* Spice Code nodes in cell cell 'inv{sch}'
#.INCLUDE Modelos_Transistores.txt
#.PARAM SUPPLY=5v
#VDD VDD 0 DC 'SUPPLY'
#Vin Vin 0 PULSE 0 'SUPPLY' 100MS 10MS 10MS 200MS 500MS
#.TRAN 1MS 600MS
.ENDS ADCD_Hipperdinger__inv

*** SUBCIRCUIT ADCD_Hipperdinger__Delayer FROM CELL Delayer{sch}
.SUBCKT ADCD_Hipperdinger__Delayer gnd vdd Vin Vout
** GLOBAL gnd
** GLOBAL vdd
Xinv@0 gnd vdd Vin net@0 ADCD_Hipperdinger__inv
Xinv@1 gnd vdd net@0 net@6 ADCD_Hipperdinger__inv
Xinv@2 gnd vdd net@6 net@3 ADCD_Hipperdinger__inv
Xinv@3 gnd vdd net@3 net@18 ADCD_Hipperdinger__inv
Xinv@4 gnd vdd net@18 net@9 ADCD_Hipperdinger__inv
Xinv@5 gnd vdd net@9 net@15 ADCD_Hipperdinger__inv
Xinv@6 gnd vdd net@15 net@12 ADCD_Hipperdinger__inv
Xinv@7 gnd vdd net@12 Vout ADCD_Hipperdinger__inv

* Spice Code nodes in cell cell 'Delayer{sch}'
#.INCLUDE Modelos_Transistores.txt
#.PARAM SUPPLY=5v
#VDD VDD 0 DC 'SUPPLY'
#Vin Vin 0 PULSE 0 'SUPPLY' 120MS 10MS 10MS 100MS 500MS
#.TRAN 1MS 1200MS
.ENDS ADCD_Hipperdinger__Delayer

*** SUBCIRCUIT ADCD_Hipperdinger__NOR FROM CELL NOR{sch}
.SUBCKT ADCD_Hipperdinger__NOR gnd Va Vb vdd Vout
** GLOBAL gnd
** GLOBAL vdd
Mnmos-4@1 Vout Va gnd gnd NMOS L=0.6U W=1.8U
Mnmos-4@2 Vout Vb gnd gnd NMOS L=0.6U W=1.8U
Mpmos-4@0 vdd Va net@62 vdd PMOS L=0.6U W=3U
Mpmos-4@2 net@62 Vb Vout pmos-4@2_b PMOS L=0.6U W=3U

* Spice Code nodes in cell cell 'NOR{sch}'
#.INCLUDE Modelos_Transistores.txt
#.PARAM SUPPLY=5v
#VDD VDD 0 DC 'SUPPLY'
#Va Va 0 PULSE 0 'SUPPLY' 100MS 10MS 10MS 200MS 500MS
#Vb Vb 0 PULSE 0 'SUPPLY' 150MS 10MS 10MS 200MS 500MS
#.TRAN 1MS 600MS
.ENDS ADCD_Hipperdinger__NOR

*** SUBCIRCUIT ADCD_Hipperdinger__CLK_noSolp FROM CELL CLK_noSolp{sch}
.SUBCKT ADCD_Hipperdinger__CLK_noSolp C1 C2 gnd vdd Vin
** GLOBAL gnd
** GLOBAL vdd
XNOR@0 gnd net@5 C2 vdd net@17 ADCD_Hipperdinger__NOR
XNOR@1 gnd C1 net@7 vdd net@15 ADCD_Hipperdinger__NOR
Xinv@0 gnd vdd Vin net@2 ADCD_Hipperdinger__inv
Xinv@1 gnd vdd net@2 net@5 ADCD_Hipperdinger__inv
Xinv@2 gnd vdd Vin net@7 ADCD_Hipperdinger__inv
Xinv@3 gnd vdd net@17 net@9 ADCD_Hipperdinger__inv
Xinv@4 gnd vdd net@9 C1 ADCD_Hipperdinger__inv
Xinv@5 gnd vdd net@15 net@12 ADCD_Hipperdinger__inv
Xinv@6 gnd vdd net@12 C2 ADCD_Hipperdinger__inv

* Spice Code nodes in cell cell 'CLK_noSolp{sch}'
#.INCLUDE Modelos_Transistores.txt
#.PARAM SUPPLY=5v
#VDD VDD 0 DC 'SUPPLY'
#Vin Vin 0 PULSE 0 'SUPPLY' 120MS 10MS 10MS 100MS 500MS
#.TRAN 1MS 1200MS
.ENDS ADCD_Hipperdinger__CLK_noSolp

*** SUBCIRCUIT ADCD_Hipperdinger__CompPaso FROM CELL CompPaso{sch}
.SUBCKT ADCD_Hipperdinger__CompPaso gnd vdd Ven VenN Vin Vout
** GLOBAL gnd
** GLOBAL vdd
Mnmos-4@2 Vin Ven Vout gnd NMOS L=0.6U W=1.8U
Mpmos-4@2 Vout VenN Vin vdd PMOS L=0.6U W=3U
.ENDS ADCD_Hipperdinger__CompPaso

*** SUBCIRCUIT ADCD_Hipperdinger__NAND FROM CELL NAND{sch}
.SUBCKT ADCD_Hipperdinger__NAND gnd Va Vb vdd Vout
** GLOBAL gnd
** GLOBAL vdd
Mnmos-4@0 Vout Vb net@0 net@0 NMOS L=0.6U W=1.8U
Mnmos-4@1 net@0 Va gnd gnd NMOS L=0.6U W=1.8U
Mpmos-4@0 vdd Vb Vout vdd PMOS L=0.6U W=3U
Mpmos-4@1 vdd Va Vout pmos-4@1_b PMOS L=0.6U W=3U

* Spice Code nodes in cell cell 'NAND{sch}'
#.INCLUDE Modelos_Transistores.txt
#.PARAM SUPPLY=5v
#VDD VDD 0 DC 'SUPPLY'
#Va Va 0 PULSE 0 'SUPPLY' 100MS 10MS 10MS 200MS 500MS
#Vb Vb 0 PULSE 0 'SUPPLY' 150MS 10MS 10MS 200MS 500MS
#.TRAN 1MS 600MS
.ENDS ADCD_Hipperdinger__NAND

*** SUBCIRCUIT ADCD_Hipperdinger__OR_NOTANOTB FROM CELL OR_NOTANOTB{sch}
.SUBCKT ADCD_Hipperdinger__OR_NOTANOTB gnd Va Vb vdd Vout
** GLOBAL gnd
** GLOBAL vdd
XNOR@0 gnd net@2 net@0 vdd net@4 ADCD_Hipperdinger__NOR
Xinv@0 gnd vdd net@4 Vout ADCD_Hipperdinger__inv
Xinv@1 gnd vdd Va net@2 ADCD_Hipperdinger__inv
Xinv@2 gnd vdd Vb net@0 ADCD_Hipperdinger__inv
.ENDS ADCD_Hipperdinger__OR_NOTANOTB

*** SUBCIRCUIT ADCD_Hipperdinger__FFD_clrn FROM CELL FFD_clrn{sch}
.SUBCKT ADCD_Hipperdinger__FFD_clrn CLK CLRn D gnd PREn Q Qn vdd
** GLOBAL gnd
** GLOBAL vdd
XCLK_noSo@0 net@280 net@257 gnd vdd CLK ADCD_Hipperdinger__CLK_noSolp
XCompPaso@4 gnd vdd net@257 net@280 net@192 net@208 ADCD_Hipperdinger__CompPaso
XCompPaso@5 gnd vdd net@280 net@257 net@208 net@180 ADCD_Hipperdinger__CompPaso
XCompPaso@6 gnd vdd net@280 net@257 D net@198 ADCD_Hipperdinger__CompPaso
XCompPaso@7 gnd vdd net@257 net@280 net@195 net@198 ADCD_Hipperdinger__CompPaso
XNAND@0 gnd net@198 CLRn vdd net@192 ADCD_Hipperdinger__NAND
XNAND@1 gnd net@183 CLRn vdd net@180 ADCD_Hipperdinger__NAND
XOR_NOTAN@0 gnd PREn net@208 vdd net@183 ADCD_Hipperdinger__OR_NOTANOTB
XOR_NOTAN@1 gnd PREn net@192 vdd net@195 ADCD_Hipperdinger__OR_NOTANOTB
Xinv@8 gnd vdd net@180 net@174 ADCD_Hipperdinger__inv
Xinv@9 gnd vdd net@174 Qn ADCD_Hipperdinger__inv
Xinv@14 gnd vdd net@183 net@329 ADCD_Hipperdinger__inv
Xinv@15 gnd vdd net@329 Q ADCD_Hipperdinger__inv

* Spice Code nodes in cell cell 'FFD_clrn{sch}'
#.INCLUDE Modelos_Transistores.txt
#.PARAM SUPPLY=5v
#VDD VDD 0 DC 'SUPPLY'
#Vin D 0 PULSE 0 'SUPPLY' 100MS 10MS 10MS 200MS 1500MS
#Vclk CLK 0 PULSE 0 'SUPPLY' 150MS 10MS 10MS 100MS 500MS
#Vclr CLRn 0 PULSE 'SUPPLY' 0 170MS 10MS 10MS 20MS 500MS
#Vpre PREn 0 PULSE 'SUPPLY' 0 570MS 10MS 10MS 20MS 500MS
#.TRAN 1MS 1200MS
.ENDS ADCD_Hipperdinger__FFD_clrn

*** SUBCIRCUIT ADCD_Hipperdinger__XOR FROM CELL XOR{sch}
.SUBCKT ADCD_Hipperdinger__XOR gnd Va Vb vdd Vout
** GLOBAL gnd
** GLOBAL vdd
XNAND@0 gnd net@8 net@5 vdd Vout ADCD_Hipperdinger__NAND
XNAND@1 gnd Va net@0 vdd net@8 ADCD_Hipperdinger__NAND
XNAND@2 gnd net@0 Vb vdd net@5 ADCD_Hipperdinger__NAND
XNAND@3 gnd Va Vb vdd net@0 ADCD_Hipperdinger__NAND

* Spice Code nodes in cell cell 'XOR{sch}'
#.INCLUDE Modelos_Transistores.txt
#.PARAM SUPPLY=5v
#VDD VDD 0 DC 'SUPPLY'
#Va Va 0 PULSE 0 'SUPPLY' 100MS 10MS 10MS 200MS 500MS
#Vb Vb 0 PULSE 0 'SUPPLY' 150MS 10MS 10MS 200MS 500MS
#.TRAN 1MS 600MS
.ENDS ADCD_Hipperdinger__XOR

.global gnd vdd

*** TOP LEVEL CELL: 3b_counter{sch}
XDelayer@0 gnd vdd qn d ADCD_Hipperdinger__Delayer
XFFD_clrn@0 clki rst_n d gnd vdd b0 qn vdd ADCD_Hipperdinger__FFD_clrn
XFFD_clrn@1 clki rst_n net@96 gnd vdd b1 FFD_clrn@1_Qn vdd ADCD_Hipperdinger__FFD_clrn
XFFD_clrn@2 clki rst_n net@0 gnd vdd b2 FFD_clrn@2_Qn vdd ADCD_Hipperdinger__FFD_clrn
XNAND@0 gnd b0 b1 vdd net@6 ADCD_Hipperdinger__NAND
XXOR@0 gnd b0 b1 vdd net@96 ADCD_Hipperdinger__XOR
XXOR@1 gnd net@8 b2 vdd net@0 ADCD_Hipperdinger__XOR
Xinv@0 gnd vdd net@6 net@8 ADCD_Hipperdinger__inv
Xinv@1 gnd vdd CLK net@130 ADCD_Hipperdinger__inv
Xinv@2 gnd vdd net@130 clki ADCD_Hipperdinger__inv

* Spice Code nodes in cell cell '3b_counter{sch}'
.INCLUDE Modelos_Transistores.txt
.PARAM SUPPLY=5v
VDD VDD 0 DC 'SUPPLY'
Vclk CLK 0 PULSE 0 'SUPPLY' 10MS 1uS 1uS 10MS 20MS
Vclr rst_n 0 PULSE 'SUPPLY' 0 0MS 1MS 1MS 10MS 500MS
.TRAN 1MS 1200MS
.END
.END
